package facade_pkg;

  `include "types.svh"
  `include "register.svh"
  `include "reg_model.svh"
  `include "memory.svh"
  `include "dma_controller.svh"

endpackage
  
