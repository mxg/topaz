//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2022 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

parameter int unsigned ADDR_BITS=16;
parameter int unsigned INDEX_BITS=8;
parameter int unsigned SIZE = (1<<INDEX_BITS);
parameter int unsigned TAG_BITS = (ADDR_BITS - INDEX_BITS);
typedef bit [TAG_BITS-1:0] tag_t;
typedef bit[INDEX_BITS-1:0] index_t;
typedef bit [ADDR_BITS-1:0] addr_t;
parameter addr_t ADDR_MASK = 'h00000fff;

let get_index(addr_t addr) = addr & ADDR_MASK;
let get_tag(addr_t addr) = addr >> INDEX_BITS;
let make_addr(tag_t tag, index_t index, tag_t[SIZE] tags) = (tags[index] << INDEX_BITS) | index;
