//------------------------------------------------------------------------------
// FIFO protocol package
//------------------------------------------------------------------------------
package fifo_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "fifo_item.svh"
  `include "fifo_driver.svh"
  `include "fifo_monitor.svh"
  `include "fifo_talker.svh"
  `include "fifo_agent.svh"
endpackage
  
