//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2024 Mark Glasser
//
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

class reg_sequence extends uvm_sequence#(uvm_reg_item);

  `uvm_object_utils(reg_sequence)

  reg_model rm;

  function new(string name="reg_sequence");
    super.new(name);
  endfunction

  task pre_start();
    if(!uvm_resource_db#(reg_model)::read_by_name("REG", "reg_model", rm, this))
      `uvm_fatal("REG_SEQUENCE", "uanble to locate register model")
  endtask

  task body();
    bit [31:0] addr;
    bit [31:0] data;
    uvm_status_e status;
    uvm_reg_data_t value;

    addr = $urandom();
    rm.addr.write(status, addr);

    data = $urandom();
    rm.data.write(status, data);

    rm.ctrl_status.cmd.write(status, 'b01);

    rm.ctrl_status.status.read(status, value);
  endtask

endclass
