//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

class test extends uvm_component;

  `uvm_component_utils(test)

  producer p;
  consumer c;
  uvm_tlm_fifo#(packet) fifo;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    p = new("producer", this);
    c = new("consumer", this);
    fifo = new("fifo", this);
  endfunction

  function void connect_phase(uvm_phase phase);
    p.put_port.connect(fifo.blocking_put_export);
    c.get_port.connect(fifo.blocking_get_export);
  endfunction

endclass

  
