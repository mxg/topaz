
package tlm2_producer_consumer_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "initiator.svh"
  `include "target.svh"
  `include "test.svh"

endpackage
