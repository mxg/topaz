package abstract_factory_pkg;

  `include "class_family.svh"
  `include "abstract_factory.svh"
  `include "concrete_factory.svh" 

endpackage
