//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2022 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

class base_transaction;

  rand op_t op;
  rand addr_t addr;
  rand int unsigned bytes;
       byte data[];

  constraint illegal   { addr > 'hf; };
  constraint align     { (addr & 'h3) == 0; };
  constraint data_size { bytes == 8; };
  constraint address   { addr <= 'h0000ffff; };
  
  local function void post_randomize();
    if(op == READ || op == NOP)
      return;
    rand_data();
  endfunction

  local function void rand_data();
    if(bytes == 0)
      return;
    data = new [bytes];
    for(int i = 0; i < bytes; i++)
      data [i] = $urandom() & 'hff;
  endfunction

  virtual function string convert2string();
    string s;
    s = $sformatf("%08x :", addr);
    s = {s, $sformatf(" %s", op.name())};
    s = {s, $sformatf(" [%0d bytes]", bytes)};
    for(int i = 0; i < bytes; i++)
      s = {s, $sformatf(" %02x", data[i])};
    return s;
  endfunction

  virtual function void copy(base_transaction rhs);
    op    = rhs.op;
    addr  = rhs.addr;
    bytes = rhs.bytes;
    if(bytes > 0) begin
      data = new [bytes];
      for(int i = 0; i < bytes; i++)
	data[i] = rhs.data[i];
    end
  endfunction

  virtual function base_transaction clone();
    base_transaction t = new();
    t.copy(this);
  endfunction
  
endclass


  
