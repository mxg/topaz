package class_family_pkg;

  import abstract_factory_pkg::*;
  import string_factory_pkg::*;
  `include "string_factory_macros.svh"
  `include "class_family.svh"

endpackage
  
