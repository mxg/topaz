//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// cc_fsm_msi
//------------------------------------------------------------------------------
class cc_fsm_msi extends cc_fsm_base
                 implements cc_fsm_intf;

  `uvm_object_utils(cc_fsm_msi)

  function new(string name = "cc_fsm_msi");
    super.new(name);
  endfunction

  virtual function void build_state_table();

    state_table[state_M][PrRd]    = state_M;
    state_table[state_M][PrWr]    = state_M;
    state_table[state_M][BusRd]   = state_S;
    state_table[state_M][BusRdX]  = state_I;

    state_table[state_S][PrRd]    = state_S;
    state_table[state_S][PrWr]    = state_M;
    state_table[state_S][BusRd]   = state_S;
    state_table[state_S][BusUpgr] = state_I;

    state_table[state_I][PrRd]    = state_S;
    state_table[state_I][BusRd]   = state_S;
    state_table[state_I][PrWr]    = state_M;
 
  endfunction
      
endclass
