//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2021 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

virtual class abstract_class;
  pure virtual function void print();
endclass

class concrete_class_1 extends abstract_class;
  function void print();
    $display("I'm a concrete_class_1");
  endfunction
endclass

class concrete_class_2 extends abstract_class;
  function void print();
    $display("I'm a concrete_class_2");
  endfunction
endclass

class concrete_class_3 extends abstract_class;
  function void print();
    $display("I'm a concrete_class_3");
  endfunction
endclass

typedef enum{C1, C2, C3} selector_t;

function abstract_class factory(selector_t selector);
  abstract_class c;
  case(selector)
    C1: begin
      concrete_class_1 c1 = new();
      c = c1;
    end
    C2: begin
      concrete_class_2 c2 = new();
      c = c2;
    end
    C3: begin
      concrete_class_1 c3 = new();
      c = c3;
    end
  endcase
  return c;
endfunction

module top;

  initial begin
    abstract_class c;

    c = factory(C2);
    c.print();
  end
  
endmodule
