//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// packet
//
// A simple, randomizable packet
//------------------------------------------------------------------------------
class packet extends uvm_object;

  typedef enum {NOP, READ, WRITE} op_t;

  rand op_t op;
  rand bit [63:0] addr;
  rand bit [31:0] data;

  function new(string name = "packet");
    super.new(name);
  endfunction

  function string convert2string();
    return $sformatf("%5s : @%016X = %08x", op.name(), addr, data);
  endfunction

endclass

