//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// tree_visitor
//------------------------------------------------------------------------------
class tree_visitor;

  function void traverse(tree t);

    node children[$];

    if(t == null)
      return;

    visit(t);

    t.get_children(children);

    foreach(children[i]) begin
      tree t;
      $cast(t, children[i]);
      traverse(t);
    end
    
  endfunction

  function void visit(tree t);
    $display("visiting node id = %0d", t.id);
  endfunction

endclass
