//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2021 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

module top;

  import type_handle_pkg::*;
  import prototype_pkg::*;

  initial begin
    abstract_prototype p;
    populate_registry();

    p = prototype_registry::get(type_handle#(concrete_prototype_1)::get_type());
    $display("p = %s", p.convert2string());
    p = prototype_registry::get(type_handle#(concrete_prototype_2)::get_type());
    $display("p = %s", p.convert2string());
    p = prototype_registry::get(type_handle#(concrete_prototype_3)::get_type());
    $display("p = %s", p.convert2string());
  end

  function void populate_registry();
    concrete_prototype_1 c1 = new();
    concrete_prototype_2 c2 = new();
    concrete_prototype_3 c3 = new();

     c1.a = 14;
     c1.b = 22;
     c2.c = 111;
     c2.d = 88;
     c3.e = 60;
     c3.f = 90;

    prototype_registry::add(type_handle#(concrete_prototype_1)::get_type(), c1);
    prototype_registry::add(type_handle#(concrete_prototype_2)::get_type(), c2);
    prototype_registry::add(type_handle#(concrete_prototype_3)::get_type(), c3);
  endfunction
  
  
endmodule

