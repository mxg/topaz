//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// top
//------------------------------------------------------------------------------
import observer_pkg::*;

class my_subscriber extends subscriber#(string);

   local string name;
   
   function new(string nm);
      name = nm;
   endfunction

   function void update(string msg);
      $display("%s : %s", name, msg);
   endfunction

endclass

module top;

   publisher#(string) pub;
   my_subscriber sub_1;
   my_subscriber sub_2;

   initial begin
      pub = new();
      sub_1 = new("sub_1");
      sub_2 = new("sub_2");

      pub.subscribe(sub_1);
      pub.subscribe(sub_2);

      pub.notify("hi there!");
      pub.notify("so long");
   end

endmodule


   


