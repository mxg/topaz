package abstract_factory_pkg;

  `include "abstract_factory.svh"
  `include "concrete_factory.svh" 

endpackage
