//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// cc_sb_base
//------------------------------------------------------------------------------
class cc_sb_base extends uvm_subscriber#(cc_transaction);

  `uvm_component_utils(cc_sb_base)

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  virtual function void write (cc_transaction t);
  endfunction
  
endclass  

//------------------------------------------------------------------------------
// cc_sb
//------------------------------------------------------------------------------
class cc_sb#(type FSM) extends cc_sb_base;

  typedef cc_sb#(FSM) this_t;
  `uvm_component_param_utils(this_t)

  local FSM fsm;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    fsm = new();
    fsm.print_state_table();
  endfunction

  function void write (cc_transaction t);
    fsm.update_state(t.op, t.addr);
  endfunction

endclass

