package qsort_pkg;

  `include "qsort_int.svh"
  `include "qsort.svh"
  `include "qsort_comparators.svh"
  `include "qsort_test.svh" 

endpackage
