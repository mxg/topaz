class memory;

  function data_t read(addr_t addr);
  endfunction

  function write(addr_t addr, data_t data);
  endfunction
  
endclass

