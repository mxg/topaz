//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2022 Mark Glasser
//
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

class reg_driver extends uvm_component;

  uvm_seq_item_pull_port#(reg_item) seq_item_port;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    seq_item_port = new("seq_item_port", this);
  endfunction

  task run_phase(uvm_phase phase);

    reg_item item;

    forever begin
      seq_item_port.get_next_item(item);
      $display("%12t: %s", $time, item.convert2string());
      #1;
      seq_item_port.item_done();
    end
  endtask

  // function string print_item(uvm_reg_item item);
  //   string s;
  //   uvm_reg rgstr;

  //   if(!$cast(rgstr, item.element))
  //     `uvm_fatal("REG_DRIVER", "$cast failure")

  //   s = item.element_kind.name();
  //   s = {s, ": ", item.kind.name()};
  //   s = {s, " name=", item.element.get_full_name()};
  //   s = {s, $sformatf(" offset=%08x", rgstr.get_offset())};
  //   s = {s, " value={"};
  //   foreach(item.value[i]) begin
  //     s = {s, $sformatf(" %08x", item.value[i])};
  //   end
  //   s = {s, " }"};

  //   return s;
  // endfunction

endclass
