//----------------------------------------------------------------------
// FIFO sequence base
//
// Bse class for fifo sequences.  Provides convenience API for driving
// FIFO transactions.
// ----------------------------------------------------------------------
class fifo_sequence_base extends uvm_sequence#(fifo_item);

  `uvm_object_utils(fifo_sequence_base)

  function new(string name = "fifo_seq");
    super.new(name);
  endfunction

  // generate a reset transaction
  virtual task reset();
    fifo_item t = new();            // create a new item
    // populate the request transaction
    t.req_rsp = fifo_item::REQ;
    t.state = fifo_item::UNKNOWN;
    t.op = fifo_item::RST;
    t.data = '0;
    execute_transaction(t);
  endtask

  // generate a write transaction -- put a new item into the fifo.
  virtual task write(input bit[31:0] data);
    fifo_item t = new();   // create a new item
    // populate the request transaction
    t.req_rsp = fifo_item::REQ;
    t.state = fifo_item::UNKNOWN;
    t.op = fifo_item::WR;
    t.data = data;
    execute_transaction(t);
  endtask

  // generate a read transaction -- pull an item from the fifo.
  virtual task read();
    fifo_item t = new();   // create a new item
    // populate the request transaction
    t.req_rsp = fifo_item::REQ;
    t.state = fifo_item::UNKNOWN;
    t.op = fifo_item::RD;
    t.data = '0;
    execute_transaction(t);
  endtask

  // generate a no-op transaction
  virtual task nop();
    fifo_item t = new();   // create a new item
    // populate the request transaction
    t.req_rsp = fifo_item::REQ;
    t.state = fifo_item::UNKNOWN;
    t.op = fifo_item::NOP;
    t.data = '0;
    execute_transaction(t);
  endtask

  // Take care of all the details of posting a request transaction to
  // the sequencer and obtaining he response.
  task execute_transaction(fifo_item t);
    wait_for_grant();      // block until sequencer is ready for us
    send_request(t);       // hand the transaction over to the sequencer
    get_response(t);       // block until response is available
  endtask

endclass
