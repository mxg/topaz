//------------------------------------------------------------------------------
// cc_pkg
//------------------------------------------------------------------------------
package cc_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "cc_types.svh"
  `include "cc_transaction.svh"
  `include "cc_fsm_base.svh"
  `include "cc_fsm_msi.svh"
  `include "cc_fsm_mesi.svh"
  `include "cc_fsm_moesi.svh"
  `include "cc_sb.svh"
  `include "cc_env.svh"
  `include "cc_test.svh"

endpackage
  
