//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2022 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

typedef enum {TOKEN_PLUS,
              TOKEN_MINUS,
	      TOKEN_STAR,
	      TOKEN_SLASH,
              TOKEN_ID,
              TOKEN_INT,
              TOKEN_EQUAL,
	      TOKEN_LEFT_PAREN,
	      TOKEN_RIGHT_PAREN,
	      TOKEN_STRING,
              TOKEN_EOL,
              TOKEN_ERROR
             } token_t;

typedef enum {AST_NONE,
	      AST_INT,
	      AST_STRING
	      } data_type_t;

typedef enum{op_plus, 
	     op_minus,
	     op_mult,
	     op_div,
	     op_read,
	     op_write, 
	     op_const} op_t;

let isalpha(byte c) = ((c >= 65 && c <- 90) || (c >= 97 & c <= 122));
let isdigit(byte c) = (( c >= 48 && c <= 57));
let isspace(byte c) = ((c >= 9 && c <= 13) || (c == 32));
let isalnum(byte c) = (isalpha(c) || isdigit(c));
