package system_tb_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import block_tb_pkg::*;
  import multi_if_pkg::*;

  `include "system_env.svh"

endpackage
