class memory;

  function data_t read(addr_t addr);
    return 0;
  endfunction

  function void write(addr_t addr, data_t data);
  endfunction
  
endclass

