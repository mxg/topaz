//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// strategy
//------------------------------------------------------------------------------
interface class strategy;
  pure virtual function void operation();
endclass

class concrete_strategy_1 implements strategy;
  virtual function void operation();
  endfunction
endclass

class concrete_strategy_2 implements strategy;
  virtual function void operation();
  endfunction
endclass

class some_context;
  strategy stgy;
endclass

module top;

  initial begin
    concrete_strategy_1 stgy1;
    some_context ctxt;

    ctxt = new();
    stgy1 = new();
    ctxt.stgy = stgy1;

  end

endmodule

    
