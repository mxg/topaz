//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2023 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// concrete_prototype_1
//------------------------------------------------------------------------------
class concrete_prototype_1 extends abstract_prototype;

   int a;
   int b;

   function void copy(concrete_prototype_1 rhs);
      a = rhs.a;
      b = rhs.b;
   endfunction

   function abstract_prototype clone();
      concrete_prototype_1 cp = new();
      cp.copy(this);
      return cp;
   endfunction

   function string convert2string();
      return $sformatf("a = %0d  b = %0d", a, b);
   endfunction

endclass

//------------------------------------------------------------------------------
// concrete_prototype_1
//------------------------------------------------------------------------------
class concrete_prototype_2 extends abstract_prototype;

   int c;
   int d;

   function void copy(concrete_prototype_2 rhs);
      c = rhs.c;
      d = rhs.d;
   endfunction

   function abstract_prototype clone();
      concrete_prototype_2 cp = new();
      cp.copy(this);
      return cp;
   endfunction

      function string convert2string();
	 return $sformatf("c = %0d  d = %0d", c, d);
   endfunction

endclass

//------------------------------------------------------------------------------
// concrete_prototype_1
//------------------------------------------------------------------------------
class concrete_prototype_3 extends abstract_prototype;

   int e;
   int f;

   function void copy(concrete_prototype_3 rhs);
      e = rhs.e;
      f = rhs.f;
   endfunction

   function abstract_prototype clone();
      concrete_prototype_3 cp = new();
      cp.copy(this);
      return cp;
   endfunction

   function string convert2string();
      return $sformatf("e = %0d  f = %0d", e, f);
   endfunction
   
endclass
