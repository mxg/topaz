package packet_pkg;

  `include "packet.svh"
  `include "udp_pkt.svh"
  `include "tcp_pkt.svh"

endpackage
  
