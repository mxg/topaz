//------------------------------------------------------------------------------
//                 .
//               .o8
//             .o888oo  .ooooo.  oo.ooooo.   .oooo.     oooooooo
//               888   d88' `88b  888' `88b `P  )88b   d'""7d8P
//               888   888   888  888   888  .oP"888     .d8P'
//               888 . 888   888  888   888 d8(  888   .d8P'  .P
//               "888" `Y8bod8P'  888bod8P' `Y888""8o d8888888P
//                                888
//                               o888o
//
//                 T O P A Z   P A T T E R N   L I B R A R Y 
//
//    TOPAZ is a library of SystemVerilog and UVM patterns and idioms.  The
//    code is suitable for study and for copying/pasting into your own work.
//
//    Copyright 2022 Mark Glasser
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//      http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
//------------------------------------------------------------------------------

class dma_controller;

  function new();
    mem = new();
    rm = new();
  endfunction

  memory mem;
  reg_model rm;
  bit ok;

  task run();
    int unsigned bytes;
    int unsigned words;
    addr_t src_addr;
    addr_t dest_addr;
    data_t data;
    
    forever begin
      rm.interrupt.poll();
      ok = 0;
      bytes = rm.byte_count.read();
      src_addr = rm.src_addr.read();
      dest_addr = rm.dest_addr.read();

      words = bytes / 4;
      for(int i = 0; i < words; i++) begin
	data = mem.read(src_addr);
	mem.write(dest_addr, data);
	src_addr += 4;
	dest_addr += 4;
      end
      ok = 1;
    end
  endtask

  function ok_to_kill();
    return ok;
  endfunction

endclass

