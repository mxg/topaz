package class_family_pkg;

  `include "class_family.svh"

endpackage
  
