package class_family_pkg;

  import type_handle_pkg::*;
  import abstract_factory_pkg::*;
  import type_factory_pkg::*;
  `include "type_factory_macros.svh"
  `include "class_family.svh"

endpackage
  
